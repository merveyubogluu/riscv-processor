module PC_4adder(

    input wire [31:0] A,
    output wire [31:0] C

    );
    
    assign C = A + 4 ;
    
endmodule
